// ctrl_bufg.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module ctrl_bufg (
		input  wire  inclk,  //  altclkctrl_input.inclk
		output wire  outclk  // altclkctrl_output.outclk
	);

	ctrl_bufg_altclkctrl_0 altclkctrl_0 (
		.inclk  (inclk),  //  altclkctrl_input.inclk
		.outclk (outclk)  // altclkctrl_output.outclk
	);

endmodule
