// import ex_types_pkg::*;
// import connect_pkg::*;


interface tb_01_if(  input wire clk );



    task init;

    endtask
    
endinterface //tb_01_if


