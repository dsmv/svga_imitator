
package tb_01_pkg;



    // virtual     axi_stream_if   #( .bytes ( n ) )  _st0;
    // virtual     axi_stream_if   #( .bytes ( n ) )  _st1;


    int                 _cnt_wr=0;
    int                 _cnt_rd=0;
    int                 _cnt_ok=0;  
    int                 _cnt_error=0;


    task tb_01_init;
    
    endtask

    task tb_01_prepare;


    endtask


endpackage    