
module ctrl_bufg (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
